`define MYINC "test.svh"

`include `MYINC

module yo();
endmodule
