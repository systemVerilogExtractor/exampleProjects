`include "test.svh"

module adder(cin, cout, s);
endmodule
