// some comment

`include "test_common.svh"

// some other comment
