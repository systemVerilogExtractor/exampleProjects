some
tokens
here